module Instructions_memory(clock, address, instrucao);
	input clock;
	input [9:0] address;
	
	output wire [31:0] instrucao;
	integer clock0 = 0;
	reg [31:0] RAM[80:0];
	
	always @ ( posedge clock ) begin
		if (clock0==0) begin
			RAM[0] = 32'b10101000000000000000000000000000; // st 32'b101010 00000 00000 0000000000000000
			RAM[1] = 32'b10001100000000010000000000000001; // ldi 32'b100010 00000 00001 0000000000000001
			RAM[2] = 32'b00000100001000100000000000000001; // addi 32'b000001 00001 00010 0000000000000001
			RAM[3] = 32'b00000000001000100001100000001001; // mult 32'b000000 00001 00010 00011 00000 001001
			RAM[4] = 32'b00010000001000100000000000000000; // beq 32'b000100 00001 00010 0000000000000000
			RAM[5] = 32'b00011000001000100000000000000000; // bne 32'b000110 00001 00010 0000000000000000
			RAM[6] = 32'b01010000000000000000000000000010; // jump 32'b010100 00000000000000000000000010
			
			clock0 <= 0;
		end
	end
	
	assign instrucao = RAM[address];
	
endmodule