module Instructions_memory(clock, address, instrucao);
	input clock;
	input [9:0] address;
	
	output wire [31:0] instrucao;
	integer clock0 = 0;
	reg [31:0] RAM[80:0];
	
	always @ ( posedge clock ) begin
		if (clock0 == 0) begin
		// programa 1: fatorial
			RAM[0] = 32'b10101011110000000000000000000000;
			// st $30 M[0] 32'b101010 11110 00000 0000000000000000;
			RAM[1] = 32'b10001000000000000000000000000000;
			// ld $0 M[0] 32'b100010 00000 00000 0000000000000000;
			RAM[2] = 32'b10001100000000010000000000000001;
			// ldi $1, $0, 1 32'b100011 00000 00001 0000000000000001;
			RAM[3] = 32'b10001100000000100000000000000000;
			// ldi $2, $0, 0 32'b100011 00000 00010 0000000000000000;
			RAM[4] = 32'b10001100000111110000000000000001;
			// display $31, 32'b100011 00000 11111 0000000000000001;
			RAM[5] = 32'b00001000000000010000000000000010;
			// *loop sub $0, $0, $2 32'b000010 00000 00001 00000 00000 000010;
			RAM[6] = 32'b00010000000000100000000000010101;
			// beq $0 $2, fim 32'b000100 00000 00010 0000000000010101;
			RAM[7] = 32'b00000011111000011111100000000001;
			// display $31 + $1 32'b000000 11111 00001 11111 00000 000001;
			RAM[8] = 32'b00001011111000010000100000000010;
			// $1 = $31 - $1 32'b000010 11111 00001 00001 00000 000010;
			RAM[9] = 32'b01000000000000000000000000000101;
			// jump to 5 32'b010000 00000000000000000000000101;
			
		// programa 2: fibonacci
			RAM[10] = 32'b10101011110000000000000000000000;
			// st $30 M[0]   32'b101010 11110 00000 0000000000000000;
			RAM[11] = 32'b10001000000000000000000000000000;
			// ld $0 M[0]    32'b100010 00000 00000 0000000000000000;
			RAM[12] = 32'b10001100000000010000000000000001;
			// ldi $1, $0, 1 32'b100011 00000 00001 0000000000000001;
			RAM[13] = 32'b10001100000000100000000000000000;
			// ldi $2, $0, 0 32'b100011 00000 00010 0000000000000000
			RAM[14] = 32'b10001100000111110000000000000001;
			// display $31,  32'b100011 00000 11111 0000000000000001;
			RAM[15] = 32'b00001000000000010000000000000010;
			// *loop sub $0, $0, $2 32'b000010 00000 00001 00000 00000 000010;
			RAM[16] = 32'b00010000000000100000000000010101;
			// beq $0 $2, fim 32'b000100 00000 00010 0000000000010101;
			RAM[17] = 32'b00000000001000000000100000001001;
			// $1 = $1 * $0 32'b000000 00001 00000 00001 00000 001001;
			RAM[18] = 32'b10101000001000000000000000000000;
			// st $1 M[0] 32'b101010 00001 00000 0000000000000000;
			RAM[19] = 32'b10001011111000000000000000000000;
			// ld $31 M[0]    32'b100010 11111 00000 0000000000000000;
			RAM[20] = 32'b01000000000000000000000000001111;
			// jump to 15 32'b010000 00000000000000000000001111;
			
			
		// programa 3: testes
			//RAM[21] = 32'b10101000000000000000000000000000;
			// st 32'b101010 00000 00000 0000000000000000
			//RAM[22] = 32'b10001100000000010000000000000001;
			// ldi 32'b100010 00000 00001 0000000000000001
			//RAM[23] = 32'b00000100001000100000000000000001;
			// addi 32'b000001 00001 00010 0000000000000001
			//RAM[24] = 32'b00000000001000100001100000001001;
			// mult 32'b000000 00001 00010 00011 00000 001001
			//RAM[25] = 32'b00010000001000100000000000000000;
			// beq 32'b000100 00001 00010 0000000000000000
			//RAM[26] = 32'b00011000001000100000000000000000;
			// bne 32'b000110 00001 00010 0000000000000000
			//RAM[27] = 32'b01010000000000000000000000000010;
			// jump 32'b010100 00000000000000000000000010
			
			clock0 <= 0;
		end
	end
	assign instrucao = RAM[address];
endmodule