module Instructions_memory(clock, address, instrucao);
	input clock;
	input [9:0] address;
	output [31:0] instrucao;
	integer clock0 = 0;
	
	reg [31:0] RAM[80:0];
	
	always @ (posedge clock) begin
		if (clock0 == 0) begin
		// programa 1: fibonacci
			RAM[1] = 32'b100011_00000_11111_0000000000000001;
			// ldi $31, 0
			RAM[2] = 32'b101010_00000_11110_0000000000000000;
			// st user_number $30
			RAM[3] = 32'b100011_00000_11111_0000000000000001;
			// ldi display_reg $31 1
			RAM[4] = 32'b100010_00000_00000_0000000000000000;
			// ld user_number $0
			RAM[5] = 32'b100011_00000_00001_0000000000000001;
			// ldi $1, 1
			RAM[6] = 32'b100011_00000_00100_0000000000000000;
			// ldi $4, 0
			RAM[7] = 32'b100011_00000_00010_0000000000000001;
			// ldi $2, 1
			RAM[8] = 32'b100011_00000_00011_0000000000000001;
			// ldi $3, 1
			RAM[9] = 32'b000000_00000_00001_00000_00000_000010;
			// sub $0, $0, $1
			RAM[10] = 32'b000100_00000_00100_0000000000111101;
			// beq $0 $4, pqp
			RAM[11] = 32'b000000_00000_00001_00000_00000_000010;
			// sub $0, $0, $1
			RAM[12] = 32'b000100_00000_00100_0000000000111101;
			// beq $0 $4, pqp
			RAM[13] = 32'b000000_00010_00011_11111_00000_000001;
			// *loop add $31, $2, $3
			RAM[14] = 32'b000000_00000_00001_00000_00000_000010;
			// sub $0, $0, $1
			RAM[15] = 32'b000100_00000_00100_0000000000111101;
			// beq $0 $4, pqp
			RAM[16] = 32'b101010_00000_11111_0000000000000000;
			// st fibonumber $31
			RAM[17] = 32'b100010_00000_00010_0000000000000000;
			// ld fibonumber $2
			RAM[18] = 32'b000000_00010_00011_11111_00000_000001;
			// add $31, $2, $3
			RAM[19] = 32'b000000_00000_00001_00000_00000_000010;
			// sub $0, $0, $1
			RAM[20] = 32'b000100_00000_00100_0000000000111101;
			// beq $0 $4, pqp
			RAM[21] = 32'b101010_00000_11111_0000000000000000;
			// st fibonumber $31
			RAM[22] = 32'b100010_00000_00011_0000000000000000;
			// ld fibonumber $3
			RAM[23] = 32'b010000_00000000000000000000001100;
			// jump to 14
			
		// programa 2: fatorial
			RAM[25] = 32'b100011_00000_11111_0000000000000010;
			// ldi $0, 0
			RAM[26] = 32'b101010_00000_11110_0000000000000000;
			// st $30 M[0]			
			RAM[27] = 32'b100010_00000_11111_0000000000000000;
			// ld display_reg $31 user_number
			RAM[28] = 32'b100010_00000_00000_0000000000000000;
			// ld user_number $0
			RAM[29] = 32'b100011_00000_00001_0000000000000001;
			// ldi $1, 1
			RAM[30] = 32'b100011_00000_00010_0000000000000000;
			// ldi $2, 0
			RAM[31] = 32'b000000_00000_00001_00000_00000_000010;
			// *loop sub $0 = $0 - $1
			RAM[32] = 32'b000100_00000_00010_0000000000111101;
			// beq $0 $2, pqp
			RAM[33] = 32'b000000_11111_00000_11111_00000_001001;
			// $31 = $31 * $0
			RAM[34] = 32'b010000_00000000000000000000011111;
			// jump to 31
			
		// programa 3: sintetico
			RAM[35] = 32'b100011_00000_11111_0000000000000011;
			// ldi $31, 0
			RAM[36] = 32'b101010_00000_11110_0000000000000000;
			// st user_number $30 M[0]
			RAM[37] = 32'b100010_00000_11111_0000000000000000;
			//ld display_reg $31 user_number
			RAM[38] = 32'b100011_00000_00001_0000000000000010;
			// ldi $1, 2
			RAM[39] = 32'b000000_11111_00001_11111_00000_000111;
			// shift left $31 << 2
			RAM[40] = 32'b000000_11111_00001_11111_00000_001000;
			// shift left $31 >> 2
			
			clock0 <= 0;
		end
	end
	assign instrucao = RAM[address];
	
endmodule
