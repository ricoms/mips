module Instructions_memory(clock, address, instrucao);
	input clock;
	input [9:0] address;
	
	output reg [31:0] instrucao;
	//integer clock0 = 0;
	reg [31:0] RAM[80:0];
	
	always @ ( posedge clock ) begin
		if (address == 0) begin
		// programa 1: fibonacci
			RAM[0] = 32'b101010_00000_11110_0000000000000000;
			// st user_number $30 M[0] 32'b101010_00000_11110_0000000000000000;
			RAM[1] = 32'b100010_11111_11111_0000000000000000;
			// ld display_reg $31 user_number 32'b100010_11111_11111_0000000000000000;
			RAM[2] = 32'b100010_00000_00000_0000000000000000;
			// ld user_number $0 M[0] 32'b100010_00000_00000_0000000000000000;
			RAM[3] = 32'b100011_00000_00001_0000000000000001;
			// ldi $1, $0, 1 32'b100011_00000_00001_0000000000000001;
			RAM[4] = 32'b100011_00000_00010_0000000000000000;
			// ldi $2, $0, 0 32'b100011_00000_00010_0000000000000000;
			RAM[5] = 32'b000000_00000_00001_00000_00000_000010;
			// *loop sub $0, $0, $2 32'b000000_00000_00001_00000_00000_000010;
			RAM[6] = 32'b000100_00000_00010_0000000000111101;
			// beq $0 $2, fim 32'b000100_00000_00010_0000000000111101;
			RAM[7] = 32'b000000_11111_00001_11111_00000_000001;
			// sum $31 = $31 + $1 32'b000000_11111_00001_11111_00000_000001;
			RAM[8] = 32'b000000_11111_00001_00001_00000_000010;
			// sub $1 = $31 - $1 32'b000000_11111_00001_00001_00000_000010;
			RAM[9] = 32'b010000_00000000000000000000001110;
			// jump to 6 32'b010000_00000000000000000000000101;
			
		// programa 2: fatorial
			RAM[15] = 32'b101010_00000_11110_0000000000000000;
			// st $30 M[0] 32'b101010_00000_11110_0000000000000000
			RAM[16] = 32'b100010_11111_11111_0000000000000000;
			// ld display_reg $31 user_number 32'b100010_11111_11111_0000000000000000;
			RAM[17] = 32'b100010_00000_00000_0000000000000000;
			// ld user_number $0 M[0] 32'b100010_00000_00000_0000000000000000;
			RAM[18] = 32'b100011_00000_00001_0000000000000001;
			// ldi $1, $0, 1 32'b100011_00000_00001_0000000000000001;
			RAM[19] = 32'b100011_00000_00010_0000000000000000;
			// ldi $2, $0, 0 32'b100011_00000_00010_0000000000000000;
			RAM[20] = 32'b000000_00000_00001_00000_00000_000010;
			// *loop sub $0, $0, $1 32'b000000_00000_00001_00000_00000_000010;
			RAM[21] = 32'b000100_00000_00010_0000000000111101;
			// beq $0 $2, fim 32'b000100_00000_00010_0000000000111101;
			RAM[22] = 32'b000000_11111_00000_11111_00000_001001;
			// $31 = $31 * $0 32'b000000_11111_00000_11111_00000_001001;
			RAM[23] = 32'b010000_00000000000000000000001110;
			// jump to 20 32'b010000_00000000000000000000010100;
			
			
		// programa 3: sintetico
			RAM[25] = 32'b101010_00000_11110_0000000000000000;
			// st user_number $30 M[0] 32'b101010_00000_11110_0000000000000000
			RAM[22] = 32'b100010_11111_11111_0000000000000000;
			//ld display_reg $31 user_number 32'b100010_11111_11111_0000000000000000;
			RAM[23] = 32'b100011_00000_00001_0000000000000010;
			// ldi $1, $0, 2 32'b100011_00000_00001_0000000000000010;
			RAM[24] = 32'b000000_11111_00001_11111_00000_000111;
			// shift left $31 << 2  32'b000000_11111_00001_11111_00000_000111;
			RAM[25] = 32'b000000_11111_00001_11111_00000_000111;
			// shift left $31 << 2  32'b000000_11111_00001_11111_00000_001000;
			//RAM[26] = 32'b00011000001000100000000000000000;
			// bne 32'b000110 00001 00010 0000000000000000
			//RAM[27] = 32'b01010000000000000000000000000010;
			// jump 32'b010100 00000000000000000000000010
			
			//clock0 <= 0;
		end
		instrucao = RAM[address];
	end
	
endmodule
